`define LENGTH 4

package test_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh";

  `include "data.svh";
  `include "seq.svh";

  `include "scoreboard.svh";
  
  `include "driver.svh";
  `include "monitor.svh";

  `include "agent.svh";
  `include "env.svh";
  `include "test.svh";
  
  endpackage // test_pkg;